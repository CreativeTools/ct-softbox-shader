MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       0Vtcytcytcy�-�ucyo��mcyo��cy}�wcytcx>cyo��Zcyo��ucyo��ucyRichtcy        PE  L ���Q        � !
  f  �      Ŵ      �                       P         @                   @� M   t� (                            0   P�                            H� @            �                           .text   %e     f                   `.rdata  �k   �  l   j             @  @.data   �0   �     �             @  �.reloc  �   0      �             @  B                                                                                                                                                                                                                                                                                                                                                                                                        U��]�  ��������  ��������������������������U��E�� tHt	-�  3�]ù��  �����]ø   ]�U�존�U��0SV��H@�A,WR������QQ���$���   h�  �������������Au������^���Q��   ���$h�  ����������^����Q�$���   h�  �����^���Q���   j h�  ���ЉF ���Q���   j h�  ���ЉF$���Q���   j h�  ���ЉF(���Q���   j h�  ������F,���Q���   ���$h�  �����^0����Q���   ���$h�  �����^8����Q���$h�  ���   �����^@����U�E��U�P�]�h�  �Q���   �M�Q�������NH�P�VL�H�NP�P�VT�H�NX�P�U�V\�U��]��P���   �E�Ph�  �M�Q�������N`�P�Vd�H�Nh�P�Vl�H�Np�P�Vt���P���   ���$h�  �����؁h!D h�  ��ݞ�   �~)  �Fx��t>�]S���!  ��t/h!D h�  ���W)  �F|��tS����   ��t_^3�[��]� _^�����[��]� ������������ �������������U���E�E�  ���������u貜  �E�M��M�]����U���`V��~  �F���W�}��؁�������U��G�������U������U���t������܎�   �������U���ڃ~$ t����܎�   �����U��~( t����܎�   �����U��~, t������܎�   �������]���������F0�]��F@�F0�]����������ؚ  �E�������Au�������0�E�������Az
������������������������-ȁ�����������N8܎�   �E��]��E����U��E����U������]�����������Dz�5��]��������v�U��������9�  �]��E����E��)�  �E��Ё����A��   �E��E��
�  ���������u����  �E������M��m������������  �N��������Au�����/��������Az����������������������-ȁ�����������M��]���Nx���E��$P��  �G���M��$Q�N|��  � �M��U��@�M��]��@�M��]����E�����������z������F`�E��_�Fh���Fp���FH���FP���FX^��������������������M��X�M��X��]� ���U���P���H@�U�A,VWR���؁���QQ���$�B,h�  ���������Q�B,���$h�  ����� ����Q�B,���$h�  ���Ћ��Q�B0jh�  ���Ћ��Q�B0jh�  ���Ћ��Q�B0jh�  ���Ћ��Q�B0jh�  ��������Q�B,���$h�  ��������Q�B,���$h�  ����������Q�B,���$h�  ��������U��U��E��]�P�Q�RHh�  ������U��U����]��P�RH�E�Ph�  ���؁���P�B,���$h�  ������   3��E;�u�MQ��   ��_3�^��]� ��U��U�R�؁���]؉}��������]��]��]����]��r  ���U�}��}����   �I\R�E�h!D P�ы��B���   ���M�Qh�  ���ҡ����   ��U�R�Ћ��E�}��}����   �R\P�M�h!D Q�ҡ��P���   ���E�Ph�  ���ҡ����   ��U�R�ЍMQ��  ��_�   ^��]� ���������������U�존�H�A���U�VR�Ћ��Q�Jj j��E�h܂P�у�j j �U�Rhp j h'  �A  ��Ph2� ��$  ���H�A�U�R�Ѓ� ��^��]�������U��V���  �Et	V�Y  ����^]� ���������������Vjh��jh�   �|  ������t%���\  �����VH�VP���VX�V`�Vh�^p^�3�^�����������U��V�u���t���QP��Ѓ��    ^]���������̡��H��@  hﾭ���Y����������U��E��t���QP��@  �Ѓ�]����������������U�존�H���  ]��������������U�존�H��  ]�������������̡��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW� �  ������u_^]Ã} tWj V蜚  �������_�F��   ^]���U����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW�w�  ������u_^]À} tWj V��  �������_�F��   ^]����������U��M��t-�=� t�y���A�uP�(�  ��]á��P�Q�Ѓ�]��������U��E��u���MP�EPQ�$  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u0jh�j;j��������t
W���q7  �3��F��u_^]� �~ t3�9_��^]� ���H<�W�҃�3Ʌ����_�F   ^��]� �����V���F   ���H<�Q��3Ʌ����^��������������̃y t�   ËA��uË��R<P��JP�у��������U����u���H�]� ���J<�URP�A�Ѓ�]� ���������������U�졤��u���H�]Ë��J<�URP�A�Ѓ�]�U�졤��$V��u���H�1����J<�URP�A�Ѓ������Q�J�E�SP�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���[t.���B�u�HV�ы��B�P�M�Q�҃���^��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^��]���������������U�졤��$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^[��]����������������U�졤��$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^[��]��U�졤��$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h,�P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^[��]����U�존�H<�A]����������������̡��H<�Q�����V��~ u>���t���Q<P�B�Ѓ��    W�~��t����,  W�d������F    _^��������U���V�E�P���A  ��P�������M���,  ��^��]��̃=� uK����t���Q<P�B�Ѓ���    ����tV���@,  V���������    ^������������U���H���H�AS�U�V3�R�]��Ћ��Q�JSj��E�h0�P�ы��B<�P�M�Q�ҋ��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���O  �M�Q�U�R�M��(P  ���&  W�}�}���   �����   �U��ATR�Ћ�������   ���Q�J�E�P���ы��B���   ���M�Qj�U�R���Ћ��Q�J���E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Bx��W�M����E���t�E� ��t���Q�J�E�P����у���t���B�P�M�Q����҃��}� u"�E�P�M�Q�M��O  ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_���H�A�U�R�Ћ��Q�JSj��E�h0�P�ы��B<�P�M�Q�ҋ��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��N  �M�Q�U�R�M��aN  ���p  W�}��I �E����   �����   �U��ATR�Ћ�������   ���Q�J�E�P���ы��B���   ���M�Qj�U�R���Ћ��Q�J���E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Bx��W�M����E��t�E ��t���Q�J�E�P����у���t���B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�����   P�BH�Ћ��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��M  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��cL  �EP�M�Q�M�u��u�L  ����   �u���E���tA��t<��uZ�����   �M�PHQ�ҋ��Q���ȋBxV�Ѕ�u-�   ^��]Ë����   �E�JTP��VP�[�������uӍUR�E�P�M��$L  ��u�3�^��]����������V��~ u>���t���Q<P�B�Ѓ��    W�~��t���J'  W��������F    _^��������U��E��� ]�̋�� @����������@����������̅�t��j�����̡��P��  �ࡴ�P��(  ��U�존�P��   ��V�E�P�ҋuP���j&  �M��&  ��^��]� ��������̡��P��$  ��U�존�H��  ]��������������U�존�H���  ]�������������̡��H��  ��U�존�H���  ]��������������U�존�H��x  ]��������������U�존�H��|  ]�������������̡��H��d  ��U�존�H��p  ]��������������U�존�H��t  ]��������������U���EV���@�t	V��������^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���I  �����   �ESP�M��#  ���Q�J�E�P�ы��B�Pj j��M�hp�Q�҃��E�P�M��l#  j j��M�Q�U�R��d���P��8  ��P�M�Q��'  ��P�U�R�'  ���P�J  ���M����#  �M��#  ��d����#  �M��#  ���H�A�U�R�Ѓ��M��j#  ��[t	V�H  ����^��]� ���U��EVP���aS  �����^]� �����Q�H  Y���������U��E�M�U�H4�M�P �U��M�@- �@8`2 �@<�2 �@@�2 �@D 2 �@H�2 �@Lp2 �@P02 �@l�2 �@X 3 �@\@2 �@`�2 �@d�2 �@T�2 �@h�2 �@p2 �@tP2 �P0�H(�@,    ]��������������U���   h�   ��`���j P�ă  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�e`  ��8��]��������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������h�Ph D �x  ���������������Vh�h�   h D ���ix  ����t���   ��t��^��3�^����������������Vh�h�   h D ���)x  ����t���   ��t��^��3�^����������������Vh�h�   h D ����w  ����t���   ��t��^��^��U��Vh�h�   h D ���w  ����t���   ��t�MQ����^]� 3�^]� �Vh�h�   h D ���yw  ����t���   ��t��^��^��U���Vh�h�   h D ���Cw  ����tI���   ��t?�E���M��$Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� ��E�^�P�X��]� ���������������Vh�h�   h D ���v  ����t���   ��t��^��3�^����������������Vh�h�   h D ���yv  ����t���   ��t��^��3�^����������������U��Vh�h�   h D ���6v  ����t���   ��t�MQ����^]� ���^]� U��Vh�h�   h D ����u  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   h D ���u  ����t���   ��t�MQ����^]� 3�^]� �U���8Vh�h�   h D ���su  ����t-���   ��t#�MWQ�U�R���Ћ��E�   ���_^��]� �E����@0    �P^�P������������X�X�X�X �؁�X(��]� ���U��Vh�h�   h D ����t  ����t���   ��t�M�UQR����^]� ����U���Vh�h�   h D ���t  ����t[���   ��tQ�MQ�U�R���Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у���^��]� �E�     �@    ^��]� ����������U��Vh�h�   h D ���t  ����t���   ��t�M�UQR����^]� 3�^]� �������������Vh�h�   h D ���s  ����t���   ��t��^��3�^����������������Vh�h�   h D ���ys  ����t���   ��t��^��3�^����������������h�h�   h D �<s  ����t���   ��t��3��������U��h�h�   h D �	s  ����t���   ��t V�u�Q�Ѓ��    ^]ËU�    ]ËE�     ]��������������Vh�h�   h D ���r  ����t���   ��t��^��3�^����������������Vh�h�   h D ���ir  ����t���   ��t��^��^��U��E�MVh!D P�  ����t+h�h�   h D �!r  ����t���   ��t��^]��^]��������Vh�h�   h D ����q  ����t���   ��t��^��3�^����������������U��Vh�h�   h D ���q  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   h D ���fq  ����t���   ��t�MQ����^]� ���^]� U��Vh�h�   h D ���&q  ����t���   ��t�M�UQR����^]� ���̡��P�BVj j����Ћ�^���������U�존�P�E�RVj P���ҋ�^]� U�존�P�E�RVPj����ҋ�^]� ���P�B�����U�존�P���   Vj ��Mj V�Ћ�^]� �����������U�존�P�EPQ�J�у�]� ����U�존�P�EPQ�J�у����@]� ���������������U�존�P�E�RtP�ҋ����   P�BX�Ѓ�]� ���U�존�P�E�Rlh#  P�EP��]� ���������������U�존�P�E�RlhF  P�EP��]� ���������������U�존�P�E�RtP�ҋ����   �M�R`QP�҃�]� ���������������U�존�P���   ]��������������U�존�P�E���   P�҅�u]� �����   P�B�Ѓ�]� ��������3�� �����������3�� ������������ �������������U����E��P�X]� �����������̸   � ��������3�� �����������3�� ������������ �������������� �������������3�� �����������U��E�M�UV�uP�EQj RPV�Q�����ǆ�   �> ǆ�   ? ǆ�   �> ǆ�   �> ǆ�   �> ǆ�    ? ǆ�   �> ǆ�   0? ǆ�   �> ǆ�    ? ^]��������U�존�P�B<��   V�uW���Ћ}��tj VW��������u_^��]�h   ������j Q�#w  �U �E�MR�UPQR������P�����Uh   ������QRWj��S  ��4_^��]������̋�`L����������̋�`\����������̋�`P����������̋�``����������̋�`D����������̋�`T����������̋�`d����������̋�`H����������̋�`X����������̋�`h���������������������������h�PhD �Pl  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�jhD �|k  ����t
�@��t]��3�]��������Vh�j\hD ���Lk  ����t�@\��tV�Ѓ���^�����Vh�j`hD ���k  ����t�@`��tV�Ѓ�^�������U��Vh�jdhD ����j  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�jhhD ���j  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�jlhD ���lj  ����t�@l��tV�Ѓ�^�������U��Vh�h�   hD ���6j  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h�   hD ����i  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�jphD ���i  ����t�@p��t�MQV�Ѓ�^]� ��^]� ��U��Vh�jxhD ���Yi  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�j|hD ���i  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�j|hD ����h  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh�h�   hD ���h  ����t=���   ��t3�MQ�U�VR��h�j`hD �Vh  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h�jhD �h  ����t	�@��t��3��������������U��V�u�> t+h�jhD ��g  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�jhD �g  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�jhD ���Ig  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�jhD ���	g  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�j hD ����f  ����t�@ ��tV�Ѓ�^�3�^���Vh�j$hD ���f  ����t�@$��tV�Ѓ�^�3�^���U��Vh�j(hD ���if  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j,hD ���f  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�j(hD ����e  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�j4hD ���e  ����t�@4��tV�Ѓ�^�3�^���U��Vh�j8hD ���Ye  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�j<hD ���	e  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�jDhD ����d  ����t�@D��tV�Ѓ�^�3�^���U��Vh�jHhD ���d  ����t�M�PHQV�҃�^]� U��Vh�jLhD ���id  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�jPhD ���)d  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�jThD ����c  ����u^Ë@TV�Ѓ�^���������U��Vh�jXhD ���c  ����t�M�PXQV�҃�^]� U��Vh�h�   hD ���c  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�h�   hD ���6c  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�h�   hD ����b  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���b  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���fb  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���&b  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�h�   hD ��a  ����u���H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]��U��Vh�h�   hD ���Va  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���a  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ����`  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���`  ����t���   ��t�MQ����^]� 3�^]� �Vh�h�   hD ���I`  ����t���   ��t��^��3�^����������������U��Vh�h�   hD ���`  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���_  ����t���   ��t�MQ����^]� ��������U��Vh�h�   hD ���v_  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�h�   hD ���)_  ����t���   ��t��^��3�^����������������VW��3����$    �h�jphD ��^  ����t�@p��t	VW�Ѓ�����8 tF��_��^�������U��SW��3�V��    h�jphD �^  ����t�@p��t	WS�Ѓ�����8 tqh�jphD �]^  ����t�@p��t�MWQ�Ѓ������h�jphD �+^  ����t�@p��t	WS�Ѓ����V���������tG�]����E^��t�8��~=h�jphD ��]  ����t�@p��t	WS�Ѓ�����8 u_�   []� _3�[]� ����������U��Vh�j\hD ���]  ����t3�@\��t,V��h�jxhD �g]  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�j\hD ���)]  ����t3�@\��t,V��h�jdhD �]  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�j\hD ����\  ����tG�@\��t@V�ЋEh�jdhD �E��E�    �E�    �\  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�j\hD ���I\  ����t\�@\��tUV��h�jdhD �'\  ����t�@d��t
�MQV�Ѓ�h�jhhD ��[  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�j\hD ���[  ������   �@\��t~V��h�jdhD �[  ����t�@d��t
�MQV�Ѓ�h�jhhD �j[  ����t�@h��t
�URV�Ѓ�h�jhhD �A[  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�jthD ���[  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�j`hD ��Z  ����th�@`��ta�M�Q�Ѓ���^��]� h�j\hD �Z  �u����t4�@\��t-V��h�jdhD �xZ  ����t�@d��th�V�Ѓ���^��]� ������U���Vh�h�   hD �5Z  ����tU���   ��tK�M�UQR�M�Q�Ћu��P���h���h�j`hD ��Y  ����te�@`��t^�U�R�Ѓ���^��]�h�j\hD ��Y  �u����t3�@\��t,V��h�jxhD �Y  ����t�@x��t
�MVQ�Ѓ���^��]�����U���Vh�h�   hD ���cY  ����tR���   ��tH�MQ�U�R���ЋuP������h�j`hD �*Y  ����t|�@`��tu�M�Q�Ѓ���^��]� h�j\hD �E�    �E�    �E�    ��X  �u����t3�@\��t,V��h�jdhD �X  ����t�@d��t
�U�RV�Ѓ���^��]� �������������̡�V��H�QV�ҡ��H$�QDV�҃���^�����������U�존V��H�QV�ҡ��H$�QDV�ҡ��U�H$�AdRV�Ѓ���^]� ��U�존V��H�QV�ҡ��H$�QDV�ҡ��U�H$�ARV�Ѓ���^]� ��U�존V��H�QV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ѓ���^]� �̡�V��H$�QHV�ҡ��H�QV�҃�^�������������U�존�P$�EPQ�JL�у�]� ����U�존�P$�R]�����������������U�존�P$�Rl]����������������̡��P$�Bp����̡��P$�BQ�Ѓ����������������U�존�P$��VWQ�J�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]� ���U�존�P$�EPQ�J�у�]� ����U�존�P$��VWQ�J �E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U�존�P$��VWQ�J$�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o������Q$�JP�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у� _��^��]� �����̡��P$�B(Q��Yá��P$�BhQ��Y�U�존�P$�EPQ�J,�у�]� ����U�존�P$�EPQ�J0�у�]� ����U�존�P$��VWQ�Jt�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]� ���U�존�P$�EPQ�J4�у�]� ����U�존�P$�EPQ�J8�у�]� ����U�존�UV��H$�ALVR�Ѓ���^]� ��������������U�존�H�QV�uV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ћ��E�Q$�J@PV�у���^]�U�존�UV��H$�A@RV�Ѓ���^]� ��������������U�존�P$�EPQ�J<�у�]� ����U�존�P$�EPQ�J<�у����@]� ���������������U�존�P$�EP�EPQ�JP�у�]� U�존�P$�EPQ�JT�у�]� ���̡��H$�QX�����U�존�H$�A\]�����������������U�존�P$�EP�EP�EPQ�J`�у�]� �����������̡��H(�������U�존�H(�AV�u�R�Ѓ��    ^]��������������U�존�P(�R]����������������̡��P(�B�����U�존�P(�R]�����������������U�존�P(�R]�����������������U�존�P(�R ]�����������������U�존�P(�E�RjP�EP��]� ��U�존�P(�E�R$P�EP�EP��]� ���P(�B(����̡��P(�B,����̡��P(�B0�����U�존�P(�R4]�����������������U�존�P(�RX]�����������������U�존�P(�R\]�����������������U�존�P(�R`]�����������������U�존�P(�Rd]�����������������U�존�P(�Rh]�����������������U�존�P(�Rl]�����������������U�존�P(�Rx]�����������������U�존�P(���   ]��������������U�존�P(�Rt]�����������������U�존�P(�Rp]�����������������U�존�P(�BpVW�}W���Ѕ�t:���Q(�Rp�GP���҅�t"���P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U�존�P(�BtVW�}W���Ѕ�t:���Q(�Rt�GP���҅�t"���P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U�존�P(�BpSVW�}W���Ѕ���   ���Q(�Rp�GP���҅���   ���P(�Rp�GP���҅�tp���P(�Bp�_S���Ѕ�tY���Q(�Rp�CP���҅�tA���P(�Bp��S���Ѕ�t*�OQ��������t��$W��������t_^�   []� _^3�[]� ���U�존�P(�BtSVW�}W���Ѕ���   ���Q(�Rt�GP���҅���   ���P(�Rt�GP���҅�tp���P(�Bt�_S���Ѕ�tY���Q(�Rt�CP���҅�tA���P(�Bt��S���Ѕ�t*�O0Q���+�����t��HW��������t_^�   []� _^3�[]� ���U������E�    �E�    �P(�RhV�E�P���҅���   �E���uG���H�A�U�R�Ћ��Q�E�RP�M�Q�ҡ��H�A�U�R�Ѓ��   ^��]� ���Qh��hj  P���   �Ћ����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�f�����3�^��]� ���E��Q�M�j HP�EQ�JP�эU�R�4������   ^��]� �����U�존��V��H�A�U�R�Ѓ��M�Q������^��u���B�P�M�Q�҃�3���]� ���H$�E�I�U�RP�ы��B�P�M�Q�҃��   ��]� �U��Q���P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�존�P(�R8]�����������������U�존�P(�R<]�����������������U�존�P(�R@]�����������������U�존�P(�RD]�����������������U�존�P(�RH]�����������������U�존�P(�E�R|P�EP��]� ����U�존�P(�RL]�����������������U�존�P(�E���   P�EP��]� �U�존�E�P(�BT���$��]� ���U�존�E�P(�BPQ�$��]� ����̡��H(�Q�����U�존�H(�AV�u�R�Ѓ��    ^]��������������U�존�P(���   ]��������������U�존�H(�A]����������������̡��H,�Q,����̡��P,�B4�����U�존�H,�A0V�u�R�Ѓ��    ^]�������������̡��P,�B8�����U�존�P,�R<��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U�존�P,�E�R@��VWP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��̡��H,�j j �҃��������������U�존�P,�EP�EPQ�J�у�]� U�존�H,�AV�u�R�Ѓ��    ^]�������������̡��P,�B����̡��P,�B����̡��P,�B����̡��P,�B ����̡��P,�B$����̡��P,�B(�����U�존�P,�R]�����������������U�존�P,�R��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U�존�H��D  ]��������������U�존�H��H  ]��������������U�존�H��L  ]��������������U�존�H�I]�����������������U�존�H�A]�����������������U�존�H�I]�����������������U�존�H�A]�����������������U�존�H�I]�����������������U�존�H���  ]��������������U�존�H�A]�����������������U���V�u�E�P���+������Q$�J�E�P�у���u-���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�3�^��]Ë��Q�J�E�jP�у���u=�U�R��������u-���H$�AH�U�R�Ћ��Q�J�E�P�у�3�^��]Ë��B�HjV�у���u���B�HV�у����I������Q$�JH�E�P�ы��B�P�M�Q�҃��   ^��]�����������U�존�H�A ]�����������������U�존�H�I(]�����������������U�존�H��  ]��������������U�존�H��   ]��������������U�존�H��  ]��������������U�존�H��  ]��������������U�존�H�A$��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]������U�존�H���  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]���U�존�H���  ]��������������U���<��SVW�E�    ��t�E�P�   �������/���Q�J�E�P�   �ы��B$�PD�M�Q�҃��}ࡴ�H�u�QV�ҡ��H$�QDV�ҡ��H$�QLVW�҃���t)���H$�AH�U�R����Ћ��Q�J�E�P�у���t&���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�_��^[��]���U�존�H�U���  ��VWR�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]�������������̡��H���   ��U�존�H���   V�uV�҃��    ^]�������������U�존�P�]�⡴�P�B����̡��P���   ��U�존�P�R`]�����������������U�존�P�Rd]�����������������U�존�P�Rh]�����������������U�존�P�Rl]�����������������U�존�P�Rp]�����������������U�존�P�Rt]�����������������U�존�P���   ]��������������U�존�P��  ]��������������U�존�P�Rx]�����������������U�존�P���   ]��������������U�존�P�R|]�����������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P�EPQ��  �у�]� �U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U��E��t ���R P�B$Q�Ѓ���t	�   ]� 3�]� U�존�P �E�RLQ�MPQ�҃�]� U��E��u]� ���R P�B(Q�Ѓ��   ]� ������U�존�P�R]�����������������U�존�P�R]�����������������U�존�P�R]�����������������U�존�P�R]�����������������U�존�P�R]�����������������U�존�P�R]�����������������U�존�P�E�R\P�EP��]� ����U�존�P�E��  P�EP��]� �U�존�E�P�B ���$��]� ���U�존�E�P�B$Q�$��]� �����U�존�E�P�B(���$��]� ���U�존�P�R,]�����������������U�존�P�R0]�����������������U�존�P�R4]�����������������U�존�P�R8]�����������������U�존�P�R<]�����������������U�존�P�R@]�����������������U�존�P�RD]�����������������U�존�P�RH]�����������������U�존�P�RL]�����������������U�존�P�RP]�����������������U�존�P���   ]��������������U�존�P�RT]�����������������U�존�P�EPQ��  �у�]� �U�존�P���   ]��������������U�존�P���   ]��������������U�존�P�RX]����������������̡��P���   ��U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]��������������U�존�P���   ]�������������̡��P���   ��U�존�P���   ]�������������̡��P���   �ࡴ�P���   �ࡴ�P���   ��U�존�H���   ]��������������U�존�H��   ]��������������U�존�H�U�E��VWRP���  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]������������U�존�H���  ]��������������U�존�P(�BPVW�}�Q�]���E�$�Ѕ�tM���G�Q(�]�E�BPQ���$�Ѕ�t,���G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U�존�P(�BTVW�}����$���Ѕ�tE���G�Q(�BT�����$�Ѕ�t(���G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U�존�P(�BTVW�}����$���Ѕ�tr���G�Q(�BT�����$�Ѕ�tU���G�Q(�BT�����$�Ѕ�t8�OQ���������t)�W0R��������t��HW��������t_�   ^]� _3�^]� ���U�존�P(�} �R8����P��]� �U�존�P�BdS�]VW��j ���Ћ��Qh���p���   h�  V�Ћ����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ��Q(�BHV���Ѕ�t ���Q(�E�R VP���҅�t�   �3��EP袢����_��^[]� ������U�존�U�� V��H$�IWR�E�P�ы����B�P�M�Q�ҡ��H�A�U�RW�Ћ��Q�J�E�P�у��U�R����������H�A�U�R�Ѓ�_��^��]� �����������U�존���   �BXQ�Ѓ���u]� ���Q|�M�RQ�MQP�҃�]� ���U�존���   �BXQ�Ѓ���u]� ���Q|�M�R8Q�MQP�҃�]� ���U��EV��j ����Qj j P�B�ЉF����^]� ��̡�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ���Q�MP�EP�Q�JP�у��F�   ^]� ���̡��H���   ��U�존�H���   V�u�R�Ѓ��    ^]����������̡��P���   Q�Ѓ�������������U�존�P�EPQ���   �у�]� ̡��H�������U�존�H�AV�u�R�Ѓ��    ^]��������������U�존�H�AV�u�R�Ѓ��    ^]��������������U�존�P��Vh�  Q���   �E�P�ы����   �Q8P�ҋ����   ��U�R�Ѓ���^��]��������������̡��P�BQ�Ѓ����������������U�존�P�EPQ�J\�у�]� ����U�존�P�EP�EP�EP�EP�EPQ���   �у�]� �U�존�P�EP�EP�EP�EPQ�JX�у�]� �������̡��P�B Q��Y�U�존�P�EP�EP�EP�EPQ���   �у�]� �����U�존�P�EP�EP�EPQ�J�у�]� ������������U�존�H��   ]��������������U�존�P�R$]�����������������U�존�P��x  ]�������������̡��P��|  ��U�존�P�EP�EP�EP�EPQ�J(�у�]� ��������U�존�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�존�P�EP�EP�EP�EPQ�J,�у�]� ��������U�존V��H�QWV�ҍx����H�QV�ҋ��Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U�존�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�존�P�EP�EPQ�J@�у�]� U�존�P�EPQ�JD�у�]� ���̡��P�BLQ�Ѓ���������������̡��P�BLQ�Ѓ���������������̡��P�BPQ�Ѓ����������������U�존�P�EPQ�JT�у�]� ����U�존�P�EPQ�JT�у�]� ����U�존�P�EP�EPQ���   �у�]� �������������U�존�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �����   j P�BV�Ћ����   �
�E�P�у� ��^��]� ������̡��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡��H�������U�존�H�AV�u�R�Ѓ��    ^]��������������U�존�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�존�P�EPQ�J�у�]� ���̡��P�BQ��Y�U�존�P�EP�EPQ�J�у�]� U��VW���T����M�U�x@�EPQR���>����H ���_^]� �U��VW���$����M�U�xD�EPQR�������H ���_^]� �V��������xH u3�^�W�������΍xH�ܬ���H �_^�����U��V���Ŭ���xL u3�^]� W��谬���M�U�xL�EPQR��蚬���H ���_^]� �������������U��V���u����xP u���^]� W���_����M�U�xP�EP�EQRP���E����H ���_^]� ��������U��V���%����xT u���^]� W�������M�xT�EPQ��������H ���_^]� U��V�������xX u���^]� W���ϫ���xX�EP��������H ���_^]� ����U���S�]VW���t.�M��&�����菫���xL�E�P��聫���H ��ҍM��`����}��tZ���H�A�U�R�Ћ��Q�J�E�WP�ы��B�P�M�Q�҃����)����@@��t���QWP�B�Ѓ�_^[��]� ������U��V��������x` u
� }  ^]� W���ݪ���x`�EP���Ϫ���H ���_^]� ��U��VW��贪���xH�EP��親���H ���_^]� ���������U��SVW��胪���x` u� }  �#���o����x`�E���P���\����H ��ҋ����H�]�QS�҃�;�A���H�QS�҃�;�,�������M�U�xD�EPQSR�������H ���_^[]� _^�����[]� ��������������U��V���թ���xP u
�����^]� W��轩���M�U�xP�EP�EQ�MR�UPQR��蛩���H ���_^]� ��������������U��V���u����xT u
�����^]� W���]����M�xT�EPQ���K����H ���_^]� ��������������U��V���%����xX tW�������xX�EP���	����H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��)  ����t.�E�;�t'���J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡��H��   ��U�존�H��$  V�u�R�Ѓ��    ^]�����������U�존�UV��H��(  VR�Ѓ���^]� �����������U�존�P�EQ��,  P�у�]� �U�존�P�EQ��,  P�у����@]� �����������̡��H��0  �⡴�H��4  �⡴�H��p  �⡴�H��t  ��U��E��t�@�3����RP��8  Q�Ѓ�]� �����U�존�P�EPQ��<  �у�]� �U�존�P�EP�EP�EPQ��@  �у�]� ���������U�존�P�EP�EPQ��D  �у�]� �������������U�존�P�EPQ��H  �у�]� �U�존�P�E��L  ��VWPQ�M�Q�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��������������̡��P��T  Q�Ѓ�������������U�존�P�EPQ��l  �у�]� ̡��P��P  Q�Ѓ�������������U�존�P�EPQ��X  �у�]� ̡��H��\  ��U�존�H��`  V�u�R�Ѓ��    ^]�����������U�존�P�EP�EP�EP�EP�EPQ��d  �у�]� �U�존�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O������3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7��蟤���xP t$S��葤��j j �XPj�FP���}����H ���[�    �~` t���H�V`�AR�Ѓ��F`    _^������������U��SV��Fx���Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR��  ����u#���h`����H��0  h  �҃��E�~P���l����j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ���Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M��������xP u����(S���آ���UR�XP�E�Pj�NQ��������H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������jh`�h�   h�   �:�������t���,���3�����������V�������N^�������������������U��QS�]VW3��{����H�QhV�҃�����u#�H��0  h`�h�  �҃�_^3�[��]� �}�H�U�R�U�EP���   RV�Ѓ���t�9}�~#�M�<� �4�tj���F  ��t��G;}�|ݍEP������_^�   [��]� ��������������U��QS�]VW3��{����H�QhV�҃�����u#�H��0  h`�h�  �҃�_^3�[��]� �}�H�U�R�U�EP���   RV�Ѓ���tӋE;�t�3�9}�~?��E�<� t.�����QP�Bh�Ѓ���t�M�<�j���_   ��t�8F;u�|ÍUR�:�����_^�   [��]� ���������U��VW�}�7��t�������N�S���V�������    _^]�U��USV��F�����N;�~w��@�+�W������%  �yH���@u��u	�   +�����J�h�h�   ��    RP��  �ЋN����t�~_��^^��[]� _�N^[]� �^^[]� ����U�존�P8�EPQ�JD�у�]� ���̡��H8�Q<�����U�존�H8�A@V�u�R�Ѓ��    ^]�������������̡��H8�������U�존�H8�AV�u�R�Ѓ��    ^]��������������U�존�P8�EP�EP�EPQ�J�у�]� ������������U�존�P8�EP�EPQ�J�у�]� ���P8�BQ�Ѓ����������������U�존�P8�EPQ�J �у�]� ����U�존�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�존�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�존�P8�EP�EPQ�J(�у�]� U�존�P8�EP�EP�EPQ�J,�у�]� ������������U�존�P8�EP�EP�EPQ�J�у�]� ������������U�존�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�존�P8�EP�EPQ�J0�у�]� U�존�P8�EP�EP�EPQ�J4�у�]� ������������U�존�P8�EPQ�J8�у�]� ����U�존�H��x  ]��������������U�존�H��|  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H�A,]�����������������U�존�H���  ]��������������U�존�H�QV�uV�ҡ��H�Q8V�҃���^]�����̡��H�Q<�����U�존�H�I@]����������������̡��H�QD����̡��H�QH�����U�존�H�AL]�����������������U�존�H�IP]�����������������U�존�H��<  ]��������������U�존�H��,  ]��������������U�존�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡��H���   �⡴�H���  ��U�존�H�U�ER�UP�ER�UP���   Rh�6  �Ѓ�]����������������U�존�H�A]�����������������U�존�H��\  ]��������������U�존�H�AT]�����������������U�존�H�AX]�����������������U�존�H�A\]����������������̡��H�Q`�����U�존�H���  ]�������������̡��H�Qd����̡��H�Qh�����U�존�H�Al]�����������������U�존�H�Ap]�����������������U�존�H�At]�����������������U�존�H��D  ]��������������U�존�H��  ]��������������U�존�H�Ix]�����������������U�존�H��@  ]��������������U��V�u��袾�����H�U�A|VR�Ѓ���^]���������U�존�H���   ]��������������U�존�H��h  ]��������������U�존�H��d  ]��������������U�존�H���  ]�������������̡��H���   ��U�존�H��l  ]��������������U�존�H��   ]��������������U�존�H��  ]��������������U��V�u���������H���   V�҃���^]���������̡��H��`  ��U�존�H��  ]��������������U�존�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�존�H���  ]��������������U��U�E���H�E���   R���\$�E�$P�у�]�U�존�H���   ]��������������U�존�H���   ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���   ]��������������U�존�H���   ]��������������U�존�H���   ]��������������U�존�H���   ]��������������U�존�H���   ]��������������U�존�H���   ]��������������U������P�E�P�E�P�E�PQ���   �у����#E���]����������������U������P�E�P�E�P�E�PQ���   �у����#E���]����������������U������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�존�H��8  ]��������������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�존�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�존�P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ�������������U�존�P0�EP�EPQ���   �у�]� �������������U�존�P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ������������̡��H0���   ��U�존�H0���   V�u�R�Ѓ��    ^]�����������U�존�H��H  ]��������������U�존�H��T  ]�������������̡��H��p  �⡴�H���  ��U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �����   �Qj PV�ҡ����   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M�茞�����Q��X  3�VP�E�hicMCP�ы��u��u����   VP�A�U�R�Ћ����   �
�E�P�у� �M��r��������   �PT�M�Q�҃���u'�u�����������   ��U�R�Ѓ���^��]Ë����   �JT�E�P�ыu��P�����������   ��M�Q�҃���^��]���������������U�존�H��  ]��������������U�존�H��\  ]��������������U�존�H�U��t  ��V�uVR�E�P�у����3����M��k�����^��]�����U�존�H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U�존�H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�(_��^��]��U�존�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у�$��^��]���U�존�H��8  ]��������������U���  ���3ŉE��M�EPQ������h   R�R  ����x	=�  |#����H��0  h��hH  �҃��E� ���H��4  ������Rh��ЋM�3̓��  ��]�������U�존�H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U�존�H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U�존�H��p  ��4�҅���   h���M��%������P�E�R4Ph���M��ҡ��P�E�R4Ph���M��ҡ��H��X  j �U�R�E�hicMCP�ы��E�    �E�    ���   j P�A�U�R�Ћ����   �
�E�P�ы����   ��M�Q�҃�$�M�軘����]��������U�존�H��p  ��4V�҅�u���H�u�QV�҃���^��]�Wh!���M��,������P�E�R4Ph!���M��ҡ��H��X  3�V�U�R�E�hicMCP�ы��u��u����   VP�A�U�R�Ћ����   �
�E�P�ы����   �PH�M�Q�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�4�M�譗��_��^��]������U�존�H��p  ��4V�҅�u���H�u�QV�҃���^��]�Wh����M��������P�E�R4Ph����M��ҡ��H��X  3�V�U�R�E�hicMCP�ы��u��u����   VP�A�U�R�Ћ����   �
�E�P�ы����   �PH�M�Q�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�4�M�蝖��_��^��]������U�존�H��p  ��4�҅�u��]�Vh#���M��$������P�E�R4Ph#���M��ҡ��H��X  3�V�U�R�E�hicMCP�ы��u��u����   VP�A�U�R�Ћ����   �
�E�P�ы����   �P8�M�Q�ҋ����   ��U�R�Ѓ�(�M��ŕ����^��]���������������U�존�H��p  ��4�҅�u��]�Vhs���M��D������P�E�R4Phs���M��ҡ��H��X  3�V�U�R�E�hicMCP�ы��u��u����   VP�A�U�R�Ћ����   �
�E�P�ы����   �P8�M�Q�ҋ����   ��U�R�Ѓ�(�M�������^��]���������������U�존�H���  ]��������������U�존�H��@  ]��������������U�존�H���  ]��������������U��V�u���t���QP��D  �Ѓ��    ^]������U�존�H��H  ]��������������U�존�H��L  ]��������������U�존�H��P  ]��������������U�존�H��T  ]��������������U�존�H��X  ]��������������U�존�H��\  ]�������������̡��H��d  ��U�존�H��h  ]��������������U�존�H��l  ]�������������̡��H���  ��U�존�H�U���  ��VR�E�P�ыu��P���Ӓ���M�������^��]�����U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H��l  ]��������������U�존�H���  ]��������������U�존�H���  ]��������������U�존�H��$  ]��������������U�존�H��(  ]��������������U�존�H��,  ]�������������̡��H��0  �⡴�H��<  ��U�존�H���  ]�������������̡��H���  ��U�존�H���  ]������������������������������U�존�H��  ]�������������̡��H��P  ��U�존�H��`  ]�������������̡����   ���   ��Q��Y��������U�존�H�A�U��� R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�I�U�R�E�P�ы��B�P<�� �M��ҋ��Q�M�RLj�j�QP�M��ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�҃���]��������������U��E�M�UP��P�EjP������]��������������̸   �����������U��V�u��t���u6�EjP��������u3�^]Ë�������t���t��U3�;P��I#�^]�������U��EHu�E�M�����   ]� �������������U��EHV����   �$�4� �   ^]á�@����uQ�EP�w�����=�6  }�����^]Ëu��t�jh��jmj�nn������t ��耦������tV���/����   ^]���    �   ^]ËM�UQR�Xc���������H^]�^]�#c����u.�&c���z������t��� ���V�n������    �   ^]Ã��^]ÍI P� � � H� +� ˬ ����h�Ph�f �P������������������U��h�jh�f �,�������t
�@��t]�����]�������U��Vh�jh�f �����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�����E�NP�у�4�M��������^]ÍM�������^]��U��h�jh�f ��������t
�@��t]��3�]��������U��h�jh�f �\�������t
�@��t]��3�]ø� ������� ����� ����� ���]� �������� ���y� ���ۻ ���g� Ë�U�������} t�y  ��]��������������̃��$�=  �   ��ÍT$��  R��<$�D$tQf�<$t�  �   �u���=� �  �   �p��  �  �u,��� u%�|$ u���u  �"��� u�|$ u�%   �t����-`��   �=� ��  �   �p��  Z������̃=�  ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uZ�z  ��=�  t2���\$�D$%�  =�  u�<$f�$f��f���d$u�%  �����$�T$�D$�   ��ÍT$�  ��P��<$f�<$t�d  ��  ��T$��  ���   �y  ��   �  ���   �L$���S  ���  ��u���=� ��  ����   ��  �=� �|  ����   �n  ZÍT$�  �D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$��  �D$��%  ����� =  �uT$u���u���t��Q���$�\$��q�&  ��Y�a���t����  �   �B����D$%�� D$������؋D$%���D$t=�f   �l$���D$�   t�- ���t��   ���������q  ���j  �����a  ���   ��������������-`��   ���������ٱ ����u����������ٛ���u�����Ë�Q�D���&  YË�U��V��������EtV�]��Y��^]� jh���)7  �E��uz��6  ��u3��8  �+  ��u��6  ���|6  ���� ��5  ���0  ��y�'  ��� 5  ��x �2  ��xj ��-  Y��u����   �2  ��3�;�u[9=�~����}�9=@u�v/  9}u��1  �R'  �Y6  �E������   �   3�9}u�=���t�''  ��j��uY��&  h  j��+  YY��;�����V�5���5���Ѕ�tWV�'  YY� ���N��V�H  Y�������uW�n)  Y3�@�6  � jh����5  ����]3�@�E��u9���   �e� ;�t��u.�H���tWVS�ЉE�}� ��   WVS�C����E����   WVS������E��u$��u WPS����Wj S�����H���tWj S�Ѕ�t��u&WVS�������u!E�}� t�H���tWVS�ЉE��E������E���E��	PQ�)8  YYËe��E�����3��!5  Ë�U��}u�$8  �u�M�U�����Y]� ��U��S�]���woVW�=P u�c:  j�8  h�   �+  YY��t���3�@Pj �5P������u&j^9�
tS��:  Y��u���:  �0�:  �0��_^�S��:  Y�s:  �    3�[]����̋T$�L$��ti3��D$��u���   r�=� t�:  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Ë�U��} t-�uj �5P����uV��9  ����P�t9  Y�^]Ë�U��QSV�5�W�5� ���5� �؉]��֋�;���   ��+��G��ruS�:  �؍GY;�sH�   ;�s���;�rP�u��)  YY��u�C;�r>P�u���(  YY��t/��P�4����� �u�=��׉��V�ף� �E�3�_^[�Ë�Vjj �i(  YY��V���� �� ��ujX^Ã& 3�^�jh���y2  �)  �e� �u�����Y�E��E������	   �E��2  ���(  Ë�U���u���������YH]���U��WV�u�M�}�����;�v;���  ���   r�=� tWV����;�^_u�9  ��   u������r)��$�� �Ǻ   ��r����$��� �$�� ��$�t� �� 0� T� #ъ��F�G�F���G������r���$�� �I #ъ��F���G������r���$�� �#ъ���������r���$�� �I ׸ ĸ �� �� �� �� �� �� �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�� ��� �� � � �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�|� �����$�,� �I �Ǻ   ��r��+��$��� �$�|� ��� �� ܹ �F#шG��������r�����$�|� �I �F#шG�F���G������r�����$�|� ��F#шG�F�G�F���G�������V�������$�|� �I 0� 8� @� H� P� X� `� s� �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�|� ���� �� �� �� �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��;��u���M8  ��U��EV���F ��uc��   �F�Hl��Hh�N�;�t����Hpu��B  ��F;��t�F����Hpu�P;  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P�1F  ��e�F�P��D  ��Yu��P�F  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�OE  �M��E��M��H��EP��E  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�\F  @PV�V������^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M�������3�;�u"�2  j^�0��B  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�m2  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]hL�SV��E  ����ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F��_t�90uj�APQ�������}� t�E��`p�3������3�PPPPP�HA  ̋�U���,���3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0��F  ����u�)1  ��RA  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�E  ����t� ��u�E�j P�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Y���9}}�}�u;�u#�I0  j^�0�o@  �}� t�E�`p����  9}v؋E��� 9Ew	�0  j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V��3  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �E  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �[E  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���W��D  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP�C  0�F�U�����;�u��|��drj jdRP�C  0��U�F����;�u��|��
rj j
RP�qC  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�������u#��,  j^�0�=  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^��?  @PVS�����0�������} ~QV�^��?  @PVS������E����   � � ������y&�߀} u9}|�}�}������Wj0S�������}� t�E��`p�3�_^[�Ë�U���,���3ŉE��EVW�}j^V�M�Q�M�Q�p�0�A  ����u��+  �0��;  ���lS�]��u�+  �0��;  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�?  ����t� ��u�E�j VS���N�����[�M�_3�^�7����Ë�U���,���3ŉE��EV�uWj_W�M�Q�M�Q�p�0��@  ����u�+  �8�5;  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�?  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^�J����Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���������������(r�_^Ë�Vh   h   3�V�@  ����t
VVVVV�E9  ^�̀zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����t����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-`���p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR��>  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z����������������������   s��̅����������������������   v��ą�j
���� 3������U���������$�\$�   ��fD$f=p�f��fT���fs�,f�� fV�f��%�   ��%�  �Y<���f,����f(4�����  +у�ʁ�   ���  �    �� fn�f��fs����fȾ��fs�&f�� fT%p�%�   ��%�  �Y� ��Y,� ��fX4��fV%���X�fT���fs�f�� fȾ�\�f=о%�  ��%�  �Y,� ��Y� �fX4�0�fT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�fȾf���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%ȾfT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(@��Y��-��Y�f(P��X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X`�fY��\`�fY��\�����f(�`�f(5��fY�fX�fp���Y�fW���?  �X�f���X�f%��fn��YT$�Y�fs�-fp�Df(=���X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��XŃ��X��X��X�fD$�D$���fL$f��f~���fT�fs� f~Ɂ�  ���   ��� �  �� �  �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$fT$��  fn�fT��fs�4f��f�f��fv�f��%�   �� ȁ�   ��r^�� fp�f���&���f|$fd$f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=p�f���Y�f~�fs� f~��� tRfT���fT��fs�,f�� fV�%�   ��%�  �Y<���f,����f(4����> �\����Ё������ u��T$��   ��� t1��#��  ��fn�fs� f��fT$�^ʺ   �  ��#��� ��   ���fp�fW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   uefL$fT$��  fn�fT��fs�4f��f��f��fv�f��%�   =�   t#fL$f��% �  �� t������fL$f��% �  �� �G  ���fL$f��% �  �� �+  ����X��ĺ�  �  fT$f~�fs� f~ҁ����¹    �� �����fؾf��Yɺ   �H  fd$fT$fp�fW�fT�fv�f��%�   =�   ��   f~��� u fs� f~��  �?��   ��  �u���fp�fW�fT�fv�f��%�   =�   uUf��fd$% �  ��  �у� ��   �� tf��%�  =�?  r���f��%�  =�?  s�������X��º�  �cf~�fs� f~��������f���   �� t:f~�   %���=  �w%r�� w��fD$�D$���f���   ��fD$�T$�ԃ��T$���T$���$�.6  �D$��Ã� ~(=   �<  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X`����� fY��\`�fY��\�����f(�`�f(5��fY�fX�fp���Y��X��X�f%��fnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=���X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� N^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� ������fD$�D$���^�X��Y��Y��X�f��%�  �   =�  ������   �� �������fD$�D$���f�fn��Y�fs�-fV��   �����   �� tf���Y ��e���f ��Y��T���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r �ɀ� fn�fs�-��fD$�D$���fd$f�����  ���?  f��3�% �  �� �-����K�����$    ��$    �ƅp����
�u;�����ƅp����2������+  ������a���t������@u��
�t�������F  �t2��t��������x������������- �ƅp����������ݽ`������a���Au����ƅp������-*��
�uS��������
�u����������   ����
�u���u
�t���ƅp����- ���u�
�t���������������x���X��ݽ`������a���u���- �
�t���ƅp������������- �ƅp����
�u����- �������->��ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���R������ٛ���t�   ø    ���   ��V��t��V���$���$��v�   ���f���t^��t����Ë�U��QQ�EQQ�$��3  YY��uL�EQQ�$��3  �EY��Y����Dz1�EQ�؁Q�]��E��$�3  �E�Y��Y����DzjX��3�@��3��Ë�U���EV�  ���3�3��  ��9Eu:9Uuz��������z��������   ��������A�E��   ������   9Mu@9Uu;��������z�������   ������A�Eu���   ��3�F�   ��9Eu(9Uu}���U�����w����U����A�Et^�����X9MuU9UuP�EQQ�$������Y�UY������z������u!����U����Au��u���0������E���^]�jh���X  j��5  Y�e� �u�N��t/�����E��t9u,�H�JP�{���Y�v�r���Y�f �E������
   �G  Ë���j�4  Y����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����j ���� �� ��V�5���$�����u�5����V�5���(���^á�����tP�5���Ѓ���������tP�,������(3  jh ���  h|��4��u�F\��f 3�G�~�~pƆ�   CƆK  C�Fh��j�4  Y�e� �vh�0��E������>   j��3  Y�}��E�Fl��u���Fl�vl�   Y�E������   �  �3�G�uj��2  Y�j��2  YË�VW���5����������Ћ���uNh  j��  ��YY��t:V�5���5���Ѕ�tj V�����YY� ��N���	V�!���Y3�W�8�_��^Ë�V��������uj�  Y��^�jh(��  �u����   �F$��tP�����Y�F,��tP�����Y�F4��tP����Y�F<��tP����Y�F@��tP����Y�FD��tP����Y�FH��tP����Y�F\=�tP�o���Yj�2  Y�e� �~h��tW�<���u����tW�B���Y�E������W   j�G2  Y�E�   �~l��t#W��  Y;=�t��0�t�? uW�|  Y�E������   V�����Y��  � �uj�1  YËuj�1  YË�U��=���tK�} u'V�5���5$��օ�t�5���5�����ЉE^j �5���5�����u�x���������t	j P�(�]Ë�Wh|��4�����u	�����3�_�V�5@�h��W��h��W� ��h��W���h��W��փ=  �5(��t�= t�= t��u$�$���,�� A� �5�� ���������   �5P�օ���   ��  �5 �5����5� ���5����5��֣��.  ��tc�=�h� �5 ���У�����tDh  j�   ��YY��t0V�5���5���Ѕ�tj V����YY� ��N��3�@��i���3�^_Ë�U��VW3��u������Y��u'9vV�D����  ;v��������uʋ�_^]Ë�U��VW3�j �u�u�-1  ������u'9vV�D����  ;v��������uË�_^]Ë�U��VW3��u�u�e1  ��YY��u,9Et'9vV�D����  ;v��������u���_^]�̋�U��hԿ�4���thĿP�@���t�u��]Ë�U���u�����Y�u�H��j��.  Y�j��-  YË�V�������V��  V�%  V��3  V�3  V�1  V�1  ��^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=<� th<��4  Y��t
�u�<�Y�b���h(�h�����YY��uTVWhF� �d�������Y��;�s���t�Ѓ�;�r�=�  _^th� �3  Y��tj jj �� 3�]�j hP��W  j��-  Y�e� 3�@9D��   �@�E�<�} ��   �5� �5��֋؉]Ѕ�th�5� �֋��}ԉ]܉}؃��}�;�rK����9t�;�r>�7�֋��q�������5� �֋��5� ��9]�u9E�t�]܉]ЉE؋��}ԋ]���E�,��}�8�s�E� ��t�ЃE����E�<��}�@�s�E�� ��t�ЃE����E������    �} u)�D   j��+  Y�u�����} tj��+  Y��i  Ë�U��j j�u������]�jj j ������Ë�U���  �u�  Yh�   ����̋�U���LV�E�P�\�j@j ^V����YY3�;�u����  ��   ���5�;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5���@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9�}k��j@j �����YY��tQ�� ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9�|����3���~r�E�� ���t\���tW�M��	��tM��uP�X���t=����������4���E�� ��E�� �Fh�  �FP�T�����   �F�E�G�E�;�|�3ۋ���5�����t���t�N��q�F���uj�X�
�C�������P�P������tB��t>W�X���t3%�   �>��u�N@�	��u�Nh�  �FP�T���t,�F�
�N@�����C���h����5��L�3�_[^�Ã������VW�����t6��   ;�s!�p�~� tV�`����@   �N�;�r��7�����' Y����� |�_^Ã=�  u��  V�5�W3���u����   <=tGV�  Y�t���u�jGW�������YY�=$��tˋ5�S�3V�  �>=Y�Xt"jS����YY���t?VSP��  ����uG���> u��5������%� �' ��    3�Y[_^��5$������%$ �����3�PPPPP�  ̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�Q/  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�l.  Y��t��M�E�F��M��E���I.  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9� u�K  h  �HVS�L�d��� �54;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H��53�����_^[�Ë�U���SV�p���3�;�u3��wf93t��f90u���f90u�W�=l�VVV+�V��@PSVV�E��׉E�;�t8P�:���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u������Y�u�S�h��E��	S�h�3�_^[�Ë�V�p��p�W��;�s���t�Ѓ�;�r�_^Ë�V�x��x�W��;�s���t�Ѓ�;�r�_^�j h   j �t�3Ʌ����P����5P�x��%P ���h � d�5    �D$�l$�l$+�SVW���1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35��W��E� �E�   �{���t�N�38�����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���%  �E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=� t h���)  ����t�UjR�����M�U�T%  �E9Xth��W�Ӌ��V%  �E�M��H����t�N�38�����N�V�3:�o����E��H����$  �����9S�O���h��W���%  ������U��V����������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U�������e� �e� SW�N�@��  ��;�t��t	�У���eV�E�P����u�3u����3�� �3����3��E�P�|��E�3E�3�;�u�O�@����u��G  ����5���։5��^_[�Ë�U��3��M;��t
@��r�3�]Ë��]Ë�U����  ���3ŉE�SV�uWV������3�Y�����;��l  j�.+  Y���  j�+  Y��u�=���   ���   �6  hL�h  �XW�*  ������   h  ��VSf�������  ��uh�SV�O*  ����t3�PPPPP�>  V�*  @Y��<v*V�*  �E��+�j��h�+�SP�$)  ����u�h��  VW�(  ����u������VW�(  ����u�h  h��W� '  ���^SSSSS�y���j��P���;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]���  YP�����PV����M�_^3�[�j�����j�)  Y��tj�)  Y��u�=�uh�   �%���h�   ����YYË�U��E3�;�0�tA��-r�H��wjX]Ë�4�]�D���jY;��#���]�������u���Ã���s�����u���Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E��
]Ë�U���5�
����t�u��Y��t3�@]�3�]�f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U���j
����3�Ë�U��} u�����    ��  ���]��uj �5P���]�W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y������U��� �e� Wj3�Y�}��9Eu�_����    �  ����x�MV�u��t��u�;����    �`  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u��t(  ������t�M�x�E��  ��E�Pj �Z&  YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U���(  ���������5��=|f��f��f�xf�tf�%pf�-l����E ���E���E����������
  ����
��
	 ���
   �����������������������
j�i3  Yj ���h������=�
 uj�E3  Yh	 ����P������������������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�����3��ȋ��~�~�~����~���������F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ���3ŉE�SW������P�v����   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�
������C����u�j �v�������vPW������Pjj ��4  3�S�v������WPW������PW�vS�3  ��DS�v������WPW������Ph   �vS�3  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�C�����jhp������G���������Gpt�l t�wh��uj �����Y�������j�B  Y�e� �wh�u�;5��t6��tV�<���u����tV�����Y����Gh�5���u�V�0��E������   뎋u�j�  YË�U���S3�S�M����������u��   ���8]�tE�M��ap��<���u��   ����ۃ��u�E��@��   ��8]�t�E��`p���[�Ë�U��� ���3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�����   �E��0=�   r����  �t  ����  �h  ��P������V  �E�PW������7  h  �CVP�-���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u������u��+�F��t)�>����E�����D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C����Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����95��T�������M�_^3�[�:�����jh��������M���:������}�������_h�u�q����E;C�W  h   �A���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�<���u�Fh=��tP�ѻ��Y�^hS�=0����Fp��   �����   j�  Y�e� �C���C���C��3��E��}f�LCf�E�@��3��E�=  }�L����@��3��E�=   }��  ����@���5���<���u���=��tP����Y���S���E������   �0j�9  Y��%���u ����tS����Y������    ��e� �E�����Ã=�  uj��V���Y��    3�Ë�U��SV�50�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5<�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=p�th���   ;�t^9uZ���   ;�t9uP�A������   ��1  YY���   ;�t9uP� ������   �q1  YY���   �������   �����YY���   ;�tD9u@���   -�   P�ܸ�����   ��   +�P�ɸ�����   +�P軸�����   谸�������   =��t9��   uP�w-  ���   臸��YY�~P�E   ����t�;�t9uP�b���Y9_�t�G;�t9uP�K���Y���Mu�V�<���Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu��0�tV�s���Y��^�3�_]�jh����������������Fpt"�~l t�����pl��uj �[���Y�������j�  Y�e� �5���lV�Y���YY�E��E������   �j�  Y�u�Ë�U��E��]Ë�U���(  ���3ŉE�S�]W���tS�(  Y������ jL������j P誶����������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M���������������j �����������P�����u��u���tS�'  Y�M�_3�[�����Ë�Vj� �Vj�������V���P���^Ë�U���5�����t]���u�u�u�u�u�����3�PPPPP�������Ë�U����u�M�詺���E����   ~�E�Pj�u�l/  ������   �M�H���}� t�M��ap��Ë�U��=� u�E����A��]�j �u����YY]Ë�U���SV�u�M��(����]�   ;�sT�M胹�   ~�E�PjS��.  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�8/  YY��t�Ej�E��]��E� Y������ *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P��'  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=� u�E�H���w�� ]�j �u�����YY]Ë�U���(���3ŉE�SV�uW�u�}�M��ָ���E�P3�SSSSW�E�P�E�P�@9  �E�E�VP�.  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�G����Ë�U���(���3ŉE�SV�uW�u�}�M��.����E�P3�SSSSW�E�P�E�P�8  �E�E�VP�:3  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[蟷���������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��UVW��t�}��u�����j^�0�%������3�E��u����+���@��tOu��u� �����j"Y�����3�_^]Ë�U��MS�YV�u3�;�u����j^�0��������   9Ev�U�;�~��@9Ew�s���j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�v���@PWV蝲����3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0���3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f��h<  �u܉C�E��E��C�E�P�uV�������$��u�M�_�s^��3�[�´����3�PPPPP�������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�|���YË�U��E�M%����#�V�u������t$��tj j �E  YY�����j^�0�������P�u��t	��D  ����D  YY3�^]Ë�S��QQ�����U�k�l$���   ���3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����EJ  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P��I  ��h��  ��x����L  �>YYt�=�� uV��K  Y��u�6�K  Y�M�_3�^������]��[Ë�U���(3��E��E�9�t�5������T�M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �Eܔ��M��M�u�]���M��]�Q��]���Y����  �\���� "   ��  �Eܐ��M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �Eܐ���E܈��M�u��M�]���]���?  �U��E܈��W����E܄��ΉU��E܄��?����Eܔ��q�����tWItHIt9It ��t���  �E�|���E�t���Eܔ��M��u��u����Eܔ��c����E�   �������E���   �E�   �E�l��������������   �$�^�E܄���E܈���Eܐ���E�d���E�\��t����E�T��h����E�L��\����E�H���E�D���E�@��M��u�M����M�]���]�M��]�Q�E�   ��Y��u����� !   �E��^�Ð�
�
�
�
�
�
m
�
N
E
��U��QQ�E���]��E��Ë�U��f�U��  ��f#�f;�u-�EQQ�$�   HYYtHtHt3�@]�j�jX]ø   ]��M�� �  f��u�E�� u�} t����������]��E��������D��z��������@]����%���   ]Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�VW3����<�<�u��8��8h�  �0���T���tF��$|�3�@_^Ã$�8� 3����S�`�V�8�W�>��t�~tW��W�����& Y����X�|ܾ8�_���t	�~uP�Ӄ���X�|�^[Ë�U��E�4�8����]�jh���C���3�G�}�3�9Pu�����j�A���h�   ����YY�u�4�8�9t���mj�|���Y��;�u�:����    3��Pj
�X   Y�]�9u+h�  W�T���uW�!���Y�����    �]���>�W����Y�E������	   �E�������j
�)���YË�U��EV�4�8��> uP�#���Y��uj�h���Y�6���^]�����������SVW�T$�D$�L$URPQQh�d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�G  �   �C�G  �d�    ��_^[ËL$�A   �   t3�D$�H3��Ѫ��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��F  3�3�3�3�3���U��SVWj Rh�Q�,d  _^[]�U�l$RQ�t$������]� ��U��M��tj�3�X��;Es�%����    3�]��MV���uF3����wVj�5P����u2�=�
 tV�>���Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u豣��Y]�V�u��u�u谤��Y3��MW�0��uFV�uj �5P�Ȁ����u^9�
t@V����Y��t���v�V����Y�Q����    3�_^]��@�������P�����Y����(�������P�����Y�����jh������������@x��t�e� ���3�@Ëe��E������sE  ������h����dË�U��E�h�l�p�t]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5p���j h�����3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�������}؅�u����T  �h�h�U�w\���]���Y�p��Q�Ã�t2��t!Ht������    ����빾p�p��l�l�
�t�t�E�   P���E�3��}���   9E�uj�-���9E�tP����Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,����M܋����9M�}�M�k��W\�D�E����w�����E������   ��u�wdS�U�Y��]�}؃}� tj �I���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E�|]Ë�U��E��]��̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h0�h � d�    P��SVW���1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M��A����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U���$���3ŉE��ES�E��EVW�E������e� �=� �E�u}h(��̀�؅��  �=@�h�S�ׅ���   �5�P��h�S����P��h��S����P��h��S����P�֣���th��S��P�֣����M�5�;�tG9�t?P���5����֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3��;E�t)P�օ�t"�ЉE��t��;E�tP�օ�t�u��ЉE��5��օ�t�u�u��u��u����3��M�_^3�[�p����Ë�U��V�uW��t�}��u�g���j^�0������_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f�����j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�����j^�0� ������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f��K���j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u�
���j^�0�0�����_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f������j"Y���뼋�U��M��x��~��u��]á���]������    �������]Ë�U��QV�uV�3M  �E�FY��u�b���� 	   �N ����/  �@t�G���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�K  �� ;�t�K  ��@;�u�u�J  Y��uV�KJ  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�GI  ���E��M�� �F����y�M���t���t�����������������@ tjSSQ�A  #����t%�F�M��3�GW�EP�u��H  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M�������E�>�u�?*u�˰?�~����} Ճ? u�E��^�Ë�U���  ���3ŉE�S�]V�u3�W�}�u����������������������������������������������������������������������������u+�����    �3��������� t
�������`p�����7  �F@u^V�J  Y������t���t�ȃ�������������A$u����t���t�ȃ�����������@$��q���3�;��g��������������������������������
  C3�������9������y
  �B�<Xw����8����3����X�j��Y������;�� 
  �$�C'���������������������������������������������	  �� tJ��t6��t%HHt����	  �������	  �������	  �������	  �������   �	  �������	  ��*u,����������������;��l	  �������������Z	  ������k�
�ʍDЉ������?	  �������4	  ��*u&����������������;��	  ��������		  ������k�
�ʍDЉ�������  ��ItU��htD��lt��w��  ������   ��  �;luC������   �������  �������  ������ �  �<6u�{4u�������� �  �������p  <3u�{2u������������������N  <d�F  <i�>  <o�6  <u�.  <x�&  <X�  ������!�����������P��P�  Y��������Yt"�����������������C������������������������������  ��d��  �X  ��S��   tL��AtHHt$HHtHH��  �� ǅ����   �������V  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ��u�d�������������ǅ����   ��  ��X�"  HHt+���  HH��  ��������������  ������t0�G�Ph   ������P������P��G  ����tǅ����   ��G�������ǅ����   �������������|  �����������t;�H��t4������   � ������t�+���ǅ����   �7  !������,  �`�������P�M���Y�  ��p�=  �%  ��e�  ��g��   ��it|��nt.��o��  �������������ǅ����   tl������   �`�������������p��dE  ���b��������� tf������f���������ǅ����   �>  ������������@ǅ����
   �������� �  ��  ��W���  ������������@�������   ������������9�����}ǅ����   �ju��gucǅ����   �W9�����~�������������   ~=��������]  V�Ҽ��������Y��������t���������������
ǅ�����   ��5����������G�������������P��������������������P������������SP�5�����Ћ���������   t������ u������PS�5������YY������gu��u������PS�5������YY�;-u������   C������S�����ǅ����   �������*��s�n���HH�X�������  ������ǅ����'   �������ǅ����   �2���������Qƅ����0������ǅ����   ������   �������� t��������@t�G���G����G���@t��3҉�������@t��|��s����ځ�����   ������ �  ����u3�9�����}ǅ����   ���������   9�����~���������u!������u����������������t-�������RPWS�)1  ��0�������؋���9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t����u�+��������(��u�`��������������I�8 t@��u�+����������������� ��  ��������@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����+�������������u%���������������� O�0����������t���������������������������P�������2���������YYt.������u%��������������˰0O������������t��ヽ���� ������tu��~q�������������������Pj�E�P������P����A  ����u69�����t.�������������������E�P���������������� YYu��#��������������P�������������]���YY������ |2������t)�������������������� O������������t��߃����� t���������������� Y���������������t���������������r��������� t
�������`p��������M�_^3�[葓���Ð��j��7�%� Ë�U��E��t���8��  uP�r���Y]Ë�U������3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5Ԁ3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�4@  ��;�t� ��  �P訌��Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5ЀSSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�z?  ��;�th���  ���P����Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�l��E�W����Y�u������E�Y�e�_^[�M�3��a����Ë�U����u�M��[����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ���3ŉE�S3�VW�]�9]u�E� �@�E�5Ԁ3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�8>  ��;�t� ��  �P謊��Y;�t	� ��  ���؅�t��?Pj S�$�����WS�u�uj�u�օ�t�uPS�u�؀�E�S������E�Y�e�_^[�M�3��4����Ë�U����u�M��.����u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U��V�u���c  �v�����v������v�����v�����v�����v�ڊ���6�ӊ���v �ˊ���v$�Ê���v(車���v,賊���v0諊���v4裊���v蛊���v8蓊���v<苊����@�v@耊���vD�x����vH�p����vL�h����vP�`����vT�X����vX�P����v\�H����v`�@����vd�8����vh�0����vl�(����vp� ����vt�����vx�����v|������@���   ��������   �������   �������   �ى�����   �Ή�����   �É�����   踉�����   證�����   袉�����   藉�����   茉�����   聉�����   �v������   �k������   �`������   �U�����@���   �G������   �<������   �1������   �&������   �������   �������   �������   ��������   �������   �������   �و�����   �Έ�����   �È����   踈����  譈����  袈����@��  蔈����  艈����  �~�����  �s�����  �h�����   �]�����$  �R�����(  �G�����,  �<�����0  �1�����4  �&�����8  ������<  ������@  ������D  �������H  ������@��L  ������P  �և����T  �ˇ����X  �������\  赇����`  誇����^]Ë�U��V�u��tY�;p�tP臇��Y�F;t�tP�u���Y�F;x�tP�c���Y�F0;��tP�Q���Y�v4;5��tV�?���Y^]Ë�U��V�u����   �F;|�tP����Y�F;��tP����Y�F;��tP�����Y�F;��tP����Y�F;��tP�ц��Y�F ;��tP迆��Y�F$;��tP譆��Y�F8;��tP蛆��Y�F<;��tP艆��Y�F@;��tP�w���Y�FD;��tP�e���Y�FH;��tP�S���Y�vL;5��tV�A���Y^]Ë�U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�X����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M��X����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���8���3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=��O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�����+��;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5��N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3�����A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ���;����   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�����3�@�   ���e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+����M���Ɂ�   �ً��]���@u�M̋U�Y��
�� u�M̉�M�_3�[����Ë�U���8���3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=��O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�����+��;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5��N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3�����A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ���;����   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�����3�@�   ���e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+����M���Ɂ�   �ً��]���@u�M̋U�Y��
�� u�M̉�M�_3�[�q���Ë�U���|���3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u�5����    �Z���3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$�B�Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�*  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  �����`�E�;���  }�ع �E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^��x���ÍI �;D<�<�<===Q=�=�=>>�=��U���t���3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uhX��S3�PPPPP觼��3�f9U�t��   �u9Uu-hP��;�u"9UuhH��CjP�{�������u��C�h@��CjP�^�������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع����`�ۉE�f�U�u�}�M���  ��y� ��`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��o���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95���  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��s  Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�0  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�	  �EPSj �u�܀�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�9  Y����  �t�Etj�  Y����x  ����   �E��   j��  �EY�   #�tT=   t7=   t;�ub��M���� ���{L�H��M�����{,� ��2��M�����z� ����M�����z�������������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�6����M��]�� �����������}�E������S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj �   Y���3���^��[�Ë�U��}t~�}�s���� "   ]��f���� !   ]�3�Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-���]���t����-���]�������t
�-���]����t	�������؛�� t���]����jhP��g���3�9�tV�E@tH9�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%� �e��U�E�������e��U�G�����V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��SVWUj j hXV�u�Z  ]_^[��]ËL$�A   �   t2�D$�H�3��Qd��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h`Vd�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y`Vu�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ����������tj�����Y� �tjh  @j�������j�Ԋ���������U��WV�u�M�}�����;�v;���  ���   r�=� tWV����;�^_u�m�����   u������r)��$� Y�Ǻ   ��r����$�4X�$�0Y��$��X�DXpX�X#ъ��F�G�F���G������r���$� Y�I #ъ��F���G������r���$� Y�#ъ���������r���$� Y�I YY�X�X�X�X�X�X�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$� Y��0Y8YDYXY�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��Z�����$�lZ�I �Ǻ   ��r��+��$��Y�$��Z��Y�YZ�F#шG��������r�����$��Z�I �F#шG�F���G������r�����$��Z��F#шG�F�G�F���G�������V�������$��Z�I pZxZ�Z�Z�Z�Z�Z�Z�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��Z���Z�Z�Z�Z�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��QQ�EV�u�E��EWV�E��[  ���Y;�u訔��� 	   �ǋ��J�u�M�Q�u�P����E�;�u����t	P蚔��Y�ϋ�����������D0� ��E��U�_^��jhp����������]܉]��E���u�?����  �$���� 	   �Ë��   ��x;�r�����  ������ 	   �!����ы����<����������L1��t�P��  Y�e� ��D0t�u�u�u�u��������E܉U��蚓��� 	   袓���  �]܉]��E������   �E܋U��p�����u�  YË�U���  �  ���3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�-����8�����    �8�������  ������S���������L8$�����$�����?�����t��u'�M����u�ϒ���  贒���    �٢���  �D8 tjj j V������V�>  Y����  ��D���  �q~���@l3�9H�� �����P��4����3�;��`  ;�t8�?����P  ����4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P����Y��t:��4���+�M3�@;���  j��D���SP��  �������  C��@����jS��D���P�  ������n  3�PPj�M�Qj��D���QP�� ���C��@����l������=  j ��,���PV�E�P��$���� �4������
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4�������  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����/  Yf;�D����I  ��8�������� t)jXP��D����  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4������C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4������i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �l���;���   j ��(���P��+�P��5����P��$���� �4�����t�(���;�������D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48�����t��(�����D��� ��8��������D�����8��� ul��D��� t-j^9�D���u�Ռ��� 	   �݌���0�?��D�������Y�1��$���� �D@t��4����8u3��$蕌���    蝌���  ������8���+�0���[�M�_3�^�VW����jh�������]���u�a����  �F���� 	   ����   ��x;�r�:����  ����� 	   �D����ҋ����<���������D0��t�S��  Y�e� ��D0t�u�uS�n������E���ŋ��� 	   �͋���  �M���E������   �E�蠅��Ë]S�C  YË�U����h   �z��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u�8���� 	   3�]Å�x;�r����� 	   �B����ދȃ���������D��@]ø0�á�Vj^��u�   �;�}�ƣ�jP�Bz��YY����ujV�5��)z��YY����ujX^�3ҹ0������� ������|�j�^3ҹ@�W�����������������t;�t��u�1�� B����|�_3�^���
  �=< t�  �5��5P��YË�U��V�u�0�;�r"����w��+�����Q�"����N �  Y�
�� V���^]Ë�U��E��}��P������E�H �  Y]ËE�� P���]Ë�U��E�0�;�r=��w�`���+�����P�ӧ��Y]Ã� P���]Ë�U��M�E��}�`�����Q褧��Y]Ã� P���]Ë�U��E��u�.����    �S������]Ë@]á����3�9�����Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�Ĉ��j^�0�������V�u�M��S���E�9X��   f�E��   f;�v6;�t;�vWSV�N�����y���� *   �n���� 8]�t�M��ap�_^[��;�t&;�w �N���j"^�0�t���8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�l�;�t9]�j����M;�t�������z�P���;��s���;��k���WSV�RM�����[�����U��j �u�u�u�u������]��������������Q�L$+ȃ����Y�  Q�L$+ȃ����Y�  ����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����ES3�VW�E�N@  ��X�X9]�E  3ɉ]���}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�S3�;�r��s3�F�ډP��t
�U�B�U�P�M�U�E�} �X�P�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[�Ë�U��MS3�VW;�|[;�sS��������<������D0t6�<0�t0�=�u+�tItIuSj��Sj��Sj������3���o���� 	   �w�������_^[]Ë�U��E���u�[����  �@���� 	   ���]Å�x;�r�7����  ����� 	   �A����Ջ�����������Dt͋]�jh���}���}����������4���E�   3�9^u5j
����Y�]�9^uh�  �FP�T���u�]��F�E������0   9]�t������������D8P����E��b}���3ۋ}j
誡��YË�U��E�ȃ���������DP���]Ë�U��Q�=��u��  �����u���  ��j �M�Qj�MQP�����t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��M���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�Ԁ���E�u�M;��   r 8^t���   8]��f����M��ap��Z�������� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p�Ԁ���:���뺋�U��j �u�u�u�������]������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��jh���9{��3ۉ]�j蠠��Y�]�j_�}�;=�}T����9�tE���@�tP��  Y���t�E��|(������ P�`����4��-G��Y����G��E������	   �E���z���j�E���YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�z���YP�K�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV����P�A  Y��Y��3�^]�jh����y��3��}�}�j�Q���Y�}�3��u�;5���   ����98t^� �@�tVPV����YY3�B�U������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��uࡴ�4�V����YY��E������   �}�E�t�E��ny���j軝��Y�j����Y������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @h������á����t���tP���Ë�U��V�uW�����u��~���    �������D�F�t8V�����V���N  V�l���P�~  ����y�����F��tP�D���f Y�f ��_^]�jh��-x���M��3��u������u�Z~���    ���������F@t�f �E��9x���V����Y�e� V�<���Y�E��E������   �ԋuV�a���Y�jh8��w���]���u��}��� 	   ����   ��x;�r��}��� 	   ������ڋ����<���������D��t�S����Y�e� ��Dt1S�0���YP�����u���E���e� �}� t�w}���M��Z}��� 	   �M���E������   �E��=w��Ë]S�����Y�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV�Y���Y���tP����u	���   u��u�@Dtj�.���j���%���YY;�tV����YP�����u
�����3�V�u��������������Y�D0 ��tW�Y|��Y����3�_^]�jhX���u���]���u�!|���  �|��� 	   ����   ��x;�r��{���  ��{��� 	   �����ҋ����<���������D0��t�S����Y�e� ��D0tS�����Y�E���{��� 	   �M���E������   �E��pu��Ë]S����YË�U��V�u�F��t�t�v�]A���f����3�Y��F�F^]��%Ā��������h�t�B��Y����̃=� uK����t���Q<P�B�Ѓ���    ����tV��� ���V蚦������    ^�                                                                                                                                                                                                                           �� �� �� �� �� ��  � � ,� 8� F� T� ^� v� �� �� �� �� �� �� �� �� $� 2� D� \� r� �� �� �� �� �� �� � � 2� >� T� `� t� �� �� �� �� �� �� �� 
� "� :� F� T� d� t� �� �� �� �� �� �� �� � � �         �t        � <� � 3� �d        �p�e                            ���Q       w   �� ��     �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?              @      �?      �?�������?{�G�z�?       @�������?�������?333333�?��@   �. �.  / / �.  / @/ P/ 0/ �/ �/ �/ �/ `/ p/  = �< `  P 0= @= P= `= p= c:\program files\maxon\cinema 4d r14\plugins\softboxshader\source\shader\softboxshader.cpp  Xsoftbox    c:\program files\maxon\cinema 4d r14\resource\_api\c4d_resource.cpp #   M_EDITOR    ��.     �������N���������������C-DT�!	@-DT�!�?res     �������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_file.cpp �������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_misc\datastructures\basearray.h  c:\program files\maxon\cinema 4d r14\resource\_api\c4d_basebitmap.cpp   c:\program files\maxon\cinema 4d r14\resource\_api\c4d_general.h    %s         c:\program files\maxon\cinema 4d r14\resource\_api\c4d_pmain.cpp    ɮ �J�     e+000                      ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �                          �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��               ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          �� �� �� ��   K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            ��   X�	    �
   ��   `�    �   ��   `�   ��   ��   0�   ��   p�   0�   h�     �!   �x   ��y   ��z   ���   ���   ��M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     �
�
H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun       �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow  Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        0�(��������������������������������������������|�x�t�p�l�h�d�`�\�X�T�P�L�H�D�@�<�8�4�0�,�(�$� ��������������������l�L�,����������`�D�4�0�(��������������l�D����������`�4�������������GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                                                                                                                                                                                                                                                                                                ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#QNAN  1#INF   1#IND   1#SNAN  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ��`�   RSDSc'�!�H���F���   C:\Program Files\MAXON\CINEMA 4D R14\plugins\SoftboxShader\obj\softboxShader_Win32_Release.pdb             �$�@�     �       ����    @   ��        ����    @   \�           l�@�               ����$�@�    0�       ����    @   t�            L���           ������$�@�    L�       ����    @   ��            �\�            ��,�           <�D�    ��        ����    @   ,� �  � `V                     ����    ����    ����    B�     ����    ����    ������ ��     ����    ����    ����    Q�     ����    ����    ����    ��     ����    ����    ����    W� ����    f� ����    ����    ����    � ����    %� ����    ����    ����    h�     ����    ����    ����    (�     ����    ����    ����    ��     ����    ����    ����    ~�     ����    ����    ����    
    ����    ����    ������    ����    ����    ����    �    ����    ����    ����[n    ����    ����    ����ZUvU    ����    ����    ����    v\    ����    ����    ����    Fd    ����    ����    ����    �l    ����    ����    ����    �n    ����    ����    ����    xp        Dp����    ����    ����    �q    ����    ����    ����    �r    ����    ����    ����    vt��         2�  �                     �� �� �� �� �� ��  � � ,� 8� F� T� ^� v� �� �� �� �� �� �� �� �� $� 2� D� \� r� �� �� �� �� �� �� � � 2� >� T� `� t� �� �� �� �� �� �� �� 
� "� :� F� T� d� t� �� �� �� �� �� �� �� � � �     �GetCurrentThreadId  � DecodePointer �GetCommandLineA �HeapAlloc GetLastError  �HeapFree  � EncodePointer IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  EGetProcAddress  �Sleep ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime %WriteFile GetModuleFileNameW  �HeapSize  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage 9LeaveCriticalSection  � EnterCriticalSection  RtlUnwind �HeapReAlloc ?LoadLibraryW  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  �RaiseException  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll      ���Q    r�          h� l� p� 0�  ��   softboxShader.cdl c4d_main                                                                                                                    D�    .?AVNodeData@@  D�    .?AVBaseData@@  D�    .?AVShaderData@@    D�    .?AVSoftboxData@@   u�  s�  sqrt                  �?pow D�    .?AVtype_info@@             N�@���D�������������
                                                                                                   	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ���  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C   ��������������������������x�t�p�l�h�d�`�\�X�T�P�L�H�@�4�,�$�d���� �����������������	         ����������|�t�d�T�D�0�������������������������������t�h�\���P�D�4� ����������������                                                                                           ��            ��            ��            ��            ��                              p�        ��@�����0�          �      ���������              �                                                                                                                                                                                                                                                                                          P�@�.   .   h����������l��������p�������   ���5      @   �  �   ����                ��   ��   ��   ��   ��   ��!   ��   |�   t�   d�   ��   ��   H�   D�    @�   \�   T�   ��   L�   ��   ��   ��   ��   ��"   |�#   x�$   t�%   l�&   `��&         �D        � 0              �                           �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                                                                                                                                                                                                                                                                                                                               �   H0d0�0�0�0�0 11:1W1v1�1�1�122y2�2b3n3R4�4�4�4G566!6<6B6]6c6~6�6�6�6�6�67777Z7|7�7�7�7818E8h8�8�8�8�8�8 9t9�9�9�9:D:d:�:�:;�;�;�;�;C<�<�<�<=)=T=]=j=�=�=�=�=�=�=�=�=>&>E>W>r>�>�>�>�>�>??'?9?K?]?o?x?�?�?�?�?�?      $  0&080A0_0�0�0�0�0�011171I1[1m11�1�1�1�1�12$262H2Q2o2�2�2�2�2�2�23.3D3`3q3�3�3�3�3�3�3�344(4F4d4v4�4�4�4�4�4�4505F5b5t5�5�5�5�5�5 66$6-6K6l6�6�6�6�6�67!7�7�7�7�7�7�7�78!8*8=8�8�8�8�8�899D9a9�9�9�9�9:]::�:�:�:�:�:;/;f;x;<)<K<�<�<�<=!=1=D=�=�=�=�=�=>$>A>T>t>�>�?�?   0  �   0�0111%1,131:1A1H1O1V1]1d1k1r1y1�1323r3�3�3"4X4�4"5e5�5�5(6�6�6�6<7Q7�7�7"8a8�8�829|9�9�95:u:�:�:�:;$;T;t;�;�;�;<4<F<t<�<�<�=�=�=�=�=�=�=�=�=>>Q?   @  �   $0R0�0�0�021e1�1252E2�2�23J3�3�34U4�4�4555�5�56E6�6�6757u7�7�78e8�8�859u9�9�9 ::$:E:�:�:;R;�;�;%<r<�<�<=9=C=p=u=�=�=�=>9>u>�>�>�>U?y?�?�? P    060_0�0�01(1G1h1�1�1�182v2�2�2!323T3e3s3�3�3�3�3�3�34"4D4d4�4�4�4�4�4 5545T5l5�5�5�5�5�5�5 66606c6v6�6�6�6�6�6�67$7D7\7p7�7�7�7�78&848G8d8�8�8�89!949T9�9�9�9�9�9:4:T:t:�:�:�:�:�:;$;D;d;�;�;�;�;<$<><U<�<�<�<�<==5=M=d=�=�=�=>>4>�>�>�>�> ???h?�?�?�? `  (  0%0d0�0�0�0�01$1D1d1�1�1�1�12!212D2q2�2�2�2�2�2�23#313@3a3�3�3�3�3�344!444T4o4}4�4�4�4�4�4545T5t5�5�5�5�5'6@6Q6m6�6�6�6�6�6	747T7t7�7�7�7�788.8>8P8t8�8�8�8�8�8�89>9U9l9}9�9�9�9�9�9:":6:E:U:f:�:�:�:;1;D;t;�;�;�;�;�;<$<D<d<�<�<�<�<=$=D=d=�=�=�=�=>$>D>d>�>�>�>�> ?D?d?�?�?�?�? p  �   0$0D0d0�0�0�0�01$1D1d1�1�1�1�12$2D2d2�2�2�2�2�2313D3a3q3�3�3�3�3�3
44D4d4�4�4�45"5�5�5�5T6t6�6�6�6�6�647Q7d7w7�7�7�78!8O8q8�8�8�8!9D9a9t9�9�9�9:1:T:t:�:�:�:;D;d;�;�;�;�;$<T<i<x<�<�<=1=Q=q=�=�=�=>6>K>q>�>?4?t?�?�? �  �   �1�1�1 2�2�2h4�4�4�4545a5q5�5�5�5�5�5$6T6t6�6�6�6�67!7D7a7t7�7�7�8�8J9O9�9�:;%;5;�;�;�;N<=#=t=�=�=�=�=>D>a>�>�>�>?$?T?�?�?�?   �  �   0$0D0d0�0�0�0�01111D1a1q1�1�1�1�12A2Q2d2�2�2�23$3A3T3q3�3�3�3�3�3444T44�4�4�45!545T5t5�5�5�5�5D6j6�6�6�6�6747T7t7�7�7�7�778w8�8�839t9�9�9:4:a:�:�:�:�:;;$;D;d;�;�;�;�;<F<d<�<�<�<�<=4=T=t=�=�=�=�=$>B>V>f>�>�>�>�>?4?`?t?�?�?�?�? �  4  0:0m0{0�0�0�0�0�01$1>1R1b1�1�1�1�1�1$282d2|2�2�2�2�23)373F3t3�3�3�3�34 494G4V4�4�4�4�455.5d5�5�5�5�5�56D6d6�6�6�6�6747T7t7�7�7�7�7�748T8t8�8�8�8�8949T9t9�9�9�9�9�9:4:Q:d:�:�:�:�:�:�:�:;(;:;L;<<D<Q<W<�<�<�<�<==4=8=<=@=D=H=Q=t=�=>D>j>o>u>y>>�>�>�>�>�>�>�>�>�>�>�>�>�>�>0?B?�?�?�?�?�?   �  �   �0�0�0�0�12"2?2n2�2�2�2�23	33K33�3�3�3�3�34Y4�4�4)5/5>5�566$6>6E6M6�6�6�6�6�6777�7�7�7�7�7�7�7 8)8O8m8t8x8|8�8�8�8�8�8�8�8�8�8�8R9]9x99�9�9�9�9�9	::::: :$:(:,:v:|:�:�:�:�:
;;';2;�=>>�> �  |   �3�4<6B6H6�67�7,8�8�9�9::%:6:@:E:s:{:�:�:�:�:;';0;;;C;a;m;�;�;�;�;D<~<�<�<�<�<=4=T=�=n>>�>�>??D?h?q?|?�?�?   �    K0�0�01181�1�1(2g2�23+333T3�3�4�4556O6�6�6�6�67Q7�7E8�8�89(9?9_9d9<:C:O:U:a:g:p:v::�:�:�:�:�:�:�:�:�:�:�:;5;u;{;�;�;�;�;�;<<�<�<�<�<8=H=N=Z=`=p=v=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>">'>->1>7><>B>G>V>l>r>z>>�>�>�>�>�>�>�>�>�>�>�>?4?=?I?�?�?�?�?�?�? �  �    000080�0�0�0�0�0�0�0�01151@1Z1e1m1}1�1�1�1�1�122%2P2�2�2�2%3j3q3�3�3�34484\4�4�4�4�4�4
5*5O5Z5i5�5�5�5�5666�7�7�7�788s8y8�8�8	99$9)9J9O9w9�9�9�9�9�9�9:�:�:;';~;=%=2=>=F=N=Z=�=�=�=�=�=>%>/>J>R>X>f>�>�>�>�>
?V?�?�?�?�? �  �   060C0I0"1'1U1[193?3E3K3Q3W3^3e3l3s3z3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34
44&4-4�45#5�6�6�6�6�6777J7U7_7x7�7�7�7�7%888�8�89}9�9::0:B:]:e:m:�:�:�:�:�:�:�:�:;5;F;Z;�;�;=<�<T=�=�=>%>^>�>�>�?�?�?�?�?�?�?     �   |0�0�1�1�2�5�7�8�8�8�8�8X9�9�9�9�9:: :H:Q:Z:p:�:�:�:�:�:�:�:�:�:;;;^;b;f;j;n;r;v;z;~;�;�;�;�;�=�=�=�=�=�=�=>>1>E>K>T>g>�>�>???e?q?    �   |0�0�0�0_1e1q1�1�1�1222$2)2.232C2r2x2�2�2�233333#313�3�3�3)484�4�4�45!5'5 6#6.646D6I6Z6b6h6r6x6�6�6�6�6�6�6�6�6�67787:9A9G9f:m:g;
<(<N<�<�<�<�?     X   �0w2�2�23�4C7G7K7O7S7W7[7_7e7�7�7v8F9�9�9|:g>y>�>�>�>�>�>�>??/?A?S?e?w?�?�?�? 0 D   �0L1@2H2�2�3r4x455-5�5�56�6�7�7J8+9�9�9j:p:~:;1;k;�;�>�> @ 0   22222"2&2*2.22262:2G2	313A3^3�3�3�= P �   �13333I3Q3�3�4�4
505=5K5{5L6�6�657O7X7�7�78$8+83888<8@8i8�8�8�8�8�8�8�8�8�8�89 9$9(9,9�9�9�9�9�9�9�9�9:I:P:T:X:\:`:d:h:l:�:�:�:�:�:U;b;{;�;�;�;�<�<�=�=�>�>$?   ` �   �0l1<2m2�2�2�2�3�3�3X4�4�4�4�45 5-595I5P5_5k5x5�5�5�5�5�5646C6L6p6�6�6�6�7	8;*;B;b;�;�;�;<?<l<w<�<�<�<�<�<�=>^>>�>�>�>�>�>�?�?�?�? p @   J0�0�0�0�0�0j1�12(2^2h283u33�3�3�34�4�4�4�4�4�4 55   � \   1111 1$101412222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2<3@3<5@5D5   �    j?n?r?v? � 8   99$9,949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�:�: � �   @4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5   � �   �0�0111$1<1@1X1h1l1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 222$2(282<2D2\2�2�2�2�2�23$3@3L3h3�3�3�3�344(4D4H4d4h4�4�4�4�45505P5p5 � X   0000L0�0�0�0�0�0�0�0�0�0�0�0�6�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9�9�9�9�9�9�9�9�9 :::`;d;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<0=8=                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        